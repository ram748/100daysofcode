module test;


 initial begin
   if( 1'bx !== 1'b1)
      $display("True");
   //else begin
   //   $display("False");
   //end
 end


endmodule:test

